`timescale 1ns / 1ps

module instruction_memory(PC, Inst);
    input [31:0] PC;
    output reg [31:0] Inst;
    
    reg [31:0] regs[17:0];
    
    initial
        begin
    regs[0] = 32'b00000000000100000000001010010011;
    regs[1] = 32'b00000000010100101000001100110011;
    regs[2] = 32'b01000000010100110000001110110011;
    regs[3] = 32'b00000000010100111000010001100011;
    regs[4] = 32'b00000000000100101000010000010011;
    regs[5] = 32'b00000000011000101111010000110011;
    regs[6] = 32'b00000000001000101000010010010011;
    regs[7] = 32'b00000000011000101001010001100011;
    regs[8] = 32'b00000000011000101110010010110011;
    regs[9] = 32'b00000000100000000010000000100011;
    regs[10] = 32'b00000000100100000010001000100011;
    regs[11] = 32'b00000000000000000010111000000011;
    regs[12] = 32'b00000000010000000010111010000011;
        end
always @(*) begin
Inst <= regs[PC >> 2];
end
endmodule
