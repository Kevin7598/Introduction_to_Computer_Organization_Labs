`timescale 1ns / 1ps

module instruction_memory(PC, Inst);
    input [31:0] PC;
    output reg [31:0] Inst;
    
    reg [31:0] regs[80:0];
    
    initial
        begin
regs[0] <= 32'b00011001001100000000001010010011;
regs[1] <= 32'b00000000000000000000000000010011;
regs[2] <= 32'b00000000000000000000000000010011;
regs[3] <= 32'b00000000010100101000001100110011;
regs[4] <= 32'b00000000000000000000000000010011;
regs[5] <= 32'b00000000000000000000000000010011;
regs[6] <= 32'b01000000011000000000001110110011;
regs[7] <= 32'b00000000011000101111111000110011;
regs[8] <= 32'b00000000001000000000111000010011;
regs[9] <= 32'b00000000000000000000000000010011;
regs[10] <= 32'b00000000000000000000000000010011;
regs[11] <= 32'b00000001110000110001001100110011;
regs[12] <= 32'b00000000000000000000000000010011;
regs[13] <= 32'b00000000000000000000000000010011;
regs[14] <= 32'b00000000011000111110001110110011;
regs[15] <= 32'b00000000000000000000000000010011;
regs[16] <= 32'b00000000000000000000000000010011;
regs[17] <= 32'b01110011001000111111111010010011;
regs[18] <= 32'b00000000000000000000000000010011;
regs[19] <= 32'b00000000000000000000000000010011;
regs[20] <= 32'b00000000010111101101111010010011;
regs[21] <= 32'b00000000000000000000000000010011;
regs[22] <= 32'b00000000000000000000000000010011;
regs[23] <= 32'b00000001110000111101001110110011;
regs[24] <= 32'b00000000000000000000000000010011;
regs[25] <= 32'b00000000000000000000000000010011;
regs[26] <= 32'b00000001000000111001001110010011;
regs[27] <= 32'b00000000000000000000000000010011;
regs[28] <= 32'b00000000000000000000000000010011;
regs[29] <= 32'b01000001110000111101001110110011;
regs[30] <= 32'b00000000011000101001100001100011;
regs[31] <= 32'b00000000000000000000000000010011;
regs[32] <= 32'b00000000000000000000000000010011;
regs[33] <= 32'b00000000000000000000001110110011;
regs[34] <= 32'b00000010000000111000100001100011;
regs[35] <= 32'b00000000000000000000000000010011;
regs[36] <= 32'b00000000000000000000000000010011;
regs[37] <= 32'b00000011110100111101001001100011;
regs[38] <= 32'b00000000000000000000000000010011;
regs[39] <= 32'b00000000000000000000000000010011;
regs[40] <= 32'b00000000000000111000001010110011;
regs[41] <= 32'b00000000000000000000000000010011;
regs[42] <= 32'b00000000000000000000000000010011;
regs[43] <= 32'b00000001110100111100100001100011;
regs[44] <= 32'b00000000000000000000000000010011;
regs[45] <= 32'b00000000000000000000000000010011;
regs[46] <= 32'b00000000000000000000001010110011;
regs[47] <= 32'b00000000010100111001110001100011;
regs[48] <= 32'b00000000000000000000000000010011;
regs[49] <= 32'b00000000000000000000000000010011;
regs[50] <= 32'b00000000010100111000100001100011;
regs[51] <= 32'b00000000000000000000000000010011;
regs[52] <= 32'b00000000000000000000000000010011;
regs[53] <= 32'b00000000000000000000001100110011;
regs[54] <= 32'b00000001110100110100110001100011;
regs[55] <= 32'b00000000000000000000000000010011;
regs[56] <= 32'b00000000000000000000000000010011;
regs[57] <= 32'b00000001110000110101100001100011;
regs[58] <= 32'b00000000000000000000000000010011;
regs[59] <= 32'b00000000000000000000000000010011;
regs[60] <= 32'b00000000000000000000111000110011;
regs[61] <= 32'b00000000000000000000111010110011;
regs[62] <= 32'b00000001100000000000000011101111;
regs[63] <= 32'b00000000000000000000000000010011;
regs[64] <= 32'b00000000000000000000000000010011;
regs[65] <= 32'b00000010011100101000100001100011;
regs[66] <= 32'b00000000000000000000000000010011;
regs[67] <= 32'b00000000000000000000000000010011;
regs[68] <= 32'b00000000010100010010000000100011;
regs[69] <= 32'b00000000011000010000001000100011;
regs[70] <= 32'b00000000000000010010111010000011;
regs[71] <= 32'b00000000010000010000111010000011;
regs[72] <= 32'b00000000010000010100111010000011;
regs[73] <= 32'b00000000000000001000000001100111;
regs[74] <= 32'b00000000000000000000000000010011;
regs[75] <= 32'b00000000000000000000000000010011;
regs[76] <= 32'b00000000000000000000000010110011;
regs[77] <= 32'b00000000000000000000001110110011;
regs[78] <= 32'b00000000000000000000000000010011;
regs[79] <= 32'b00000000000000000000000000010011;
regs[80] <= 32'b00000000000000000000000000010011;

        end
always @(*) begin
Inst <= regs[PC >> 2];
end
endmodule
